`define ROW_A 4
`define ROW_W 4
`define COL_A 4
`define COL_W 4
`define ROW_M 16
`define COL_M 16
`define ROW_N 16
`define COL_N 16
`define EXPONENT 8
`define MANTISSA 23
`define DATA_WIDTH 16
`define WEIGHT_WIDTH 16
`define OUT_WIDTH 16
`define BUS_WIDTH 64
`define PIPELINE 0
`define DATA_TYPE 0
`define ADDR_WIDTH 32
`define A_ADDR 0
`define W_ADDR 256
`define C_ADDR 512
`define VLEN 64
`define SEW 16

